`include "JAM.v"
`include "perm_gen.sv"
