`include "SME.v"
